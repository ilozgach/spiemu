`ifndef DEFS_SVH
`define DEFS_SVH

`define ULPI_STRAP_REGISTER_ADDRESS 6'h16
`define ULPI_TX_CMD_CODE_REG_WRITE_OFFSET 8'h06
`define ULPI_TX_CMD_CODE_REG_WRITE_VALUE 2

typedef enum byte {
    ULPI_FSM_STATE_RESET,                                  // 0
    ULPI_FSM_STATE_RESET_SET_STP_HIGH,                     // 1
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_HIGH_AFTER_STP_HIGH, // 2
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_LOW_AFTER_RST_LOW,   // 3

    ULPI_FSM_STATE_WRITE_STRAP, // 4
    ULPI_FSM_STATE_READ_STRAP,  // 5

    ULPI_FSM_STATE_RX_CMD, // 6

    ULPI_FSM_STATE_REG_READ_WAIT_FOR_DIR_HIGH,   // 7
    ULPI_FSM_STATE_REG_READ_DIR_HIGH_TURNAROUND, // 8
    ULPI_FSM_STATE_REG_READ_WAIT_FOR_DIR_LOW,    // 9
    ULPI_FSM_STATE_REG_READ_DIR_LOW_TURNAROUND,  // a

    ULPI_FSM_STATE_TX_CMD_BEGIN, // b
    ULPI_FSM_STATE_TX_CMD_WAIT_NXT_HIGH, // c
    ULPI_FSM_STATE_TX_CMD_WAIT_NXT_HIGH_LAST,   // d
    ULPI_FSM_STATE_TX_CMD_END, // e

    ULPI_FSM_STATE_IDLE,               // f
    ULPI_FSM_STATE_DIR_HIGH_TURNAROUND // 10
} ulpi_fsm_state;

`endif