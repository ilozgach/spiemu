typedef enum integer {
    ULPI_FSM_STATE_RESET,
    ULPI_FSM_STATE_RESET_SET_STP_HIGH,
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_HIGH_AFTER_STP_HIGH,
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_LOW_AFTER_RST_LOW,
    ULPI_FSM_STATE_RESET_FINISH
} ulpi_fsm_state;
