typedef enum integer {
    ULPI_FSM_STATE_RESET,
    ULPI_FSM_STATE_RESET_SET_STP_HIGH,
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_HIGH_AFTER_STP_HIGH,
    ULPI_FSM_STATE_RESET_WAIT_FOR_DIR_LOW_AFTER_RST_LOW,

    ULPI_FSM_STATE_RX_CMD,

    ULPI_FSM_STATE_IDLE
} ulpi_fsm_state;
